
// 8 x 8 multiplier
module matrixMultiplier(
    input [63:0] a,
    input [63:0] b,
    output [63:0] result
);



endmodule