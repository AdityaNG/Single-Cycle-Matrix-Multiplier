
// 4 bit : 4 x 4 multiplier
module matrixMultiplier(
    input [63:0] a,
    input [63:0] b,
    output [63:0] result
);


endmodule